�]q (cpygments.token
_TokenType
qX   Keywordq�q�q�q}q(X   subtypesqcbuiltins
set
q]q	(hhX   Wordq
�q�q�q}q(hh]q�qRqX   parentqhubhhh�q�q�q}q(hh]q�qRqhhubhhX   Typeq�q�q�q}q(hh]q�q Rq!hhubhhX   PreProcq"�q#�q$�q%}q&(hh]q'�q(Rq)hhubhhX   Controlq*�q+�q,�q-}q.(hh]q/�q0Rq1hhubhhX   Constantq2�q3�q4�q5}q6(hh]q7�q8Rq9hhubhhX	   Namespaceq:�q;�q<�q=}q>(hh]q?�q@RqAhhubhhX   PseudoqB�qC�qD�qE}qF(hh]qG�qHRqIhhubhhX   DeclarationqJ�qK�qL�qM}qN(hh]qO�qPRqQhhubhhX   ReservedqR�qS�qT�qU}qV(hh]qW�qXRqYhhube�qZRq[hh)�q\�q]}q^(hh]q_(hX   Escapeq`�qa�qb�qc}qd(hh]qe�qfRqghh]ubhX   Operatorqh�qi�qj�qk}ql(hh]qm(hhhX   DBSqn�qo�qp�qq}qr(hh]qs�qtRquhhkubhhhh
�qv�qw�qx}qy(hh]qz�q{Rq|hhkube�q}Rq~hh]h
hxhnhqubhX   Nameq�q��q��q�}q�(hh]q�(hhX   Tagq��q��q��q�}q�(hh]q��q�Rq�hh�ubhhX   Entityq��q��q��q�}q�(hh]q�hhh�hn�q��q��q�}q�(hh]q��q�Rq�hh�uba�q�Rq�hh�hnh�ubhhX	   Exceptionq��q��q��q�}q�(hh]q��q�Rq�hh�ubhhX	   Decoratorq��q��q��q�}q�(hh]q��q�Rq�hh�ubhhX   Classq��q��q��q�}q�(hh]q�(hhh�hn�q��q��q�}q�(hh]q��q�Rq�hh�ubhhh�X   Startq��q��q��q�}q�(hh]q��q�Rq�hh�ube�q�Rq�hh�h�h�hnh�ubhhX   VariableqÆqąqŁq�}q�(hh]q�(hhh�X	   Anonymousqɇqʅqˁq�}q�(hh]q΅q�Rq�hh�ubhhh�h��qхqҁq�}q�(hh]qՅq�Rq�hh�ubhhh�X   Magicq؇qمqځq�}q�(hh]q݅q�Rq�hh�ubhhh�X   Globalq��q�q�q�}q�(hh]q�q�Rq�hh�ubhhh�X   Instanceq�q�q�q�}q�(hh]q�q�Rq�hh�ube�q�Rq�hh�h�h�h�h�h�h�h�h�h�h�ubhhX	   Attributeq�q�q�q�}q�(hh]q�hhh�hÇq��q��q�}q�(hh]q��q�Rq�hh�uba�q�Rr   hh�h�h�ubhhh:�r  �r  �r  }r  (hh]r  �r  Rr  hh�ubhhX   Propertyr  �r	  �r
  �r  }r  (hh]r  �r  Rr  hh�ubhhX   Symbolr  �r  �r  �r  }r  (hh]r  �r  Rr  hh�ubhhX   Classesr  �r  �r  �r  }r  (hh]r  �r  Rr  hh�ubhhhB�r   �r!  �r"  }r#  (hh]r$  �r%  Rr&  hh�ubhhX   Labelr'  �r(  �r)  �r*  }r+  (hh]r,  �r-  Rr.  hh�ubhhhh�r/  �r0  �r1  }r2  (hh]r3  �r4  Rr5  hh�ubhhX   Builtinr6  �r7  �r8  �r9  }r:  (hh]r;  (hhj6  hB�r<  �r=  �r>  }r?  (hh]r@  �rA  RrB  hj9  ubhhj6  h�rC  �rD  �rE  }rF  (hh]rG  �rH  RrI  hj9  ube�rJ  RrK  hh�hBj>  hjE  ubhhX   FieldrL  �rM  �rN  �rO  }rP  (hh]rQ  �rR  RrS  hh�ubhhX   OtherrT  �rU  �rV  �rW  }rX  (hh]rY  hhjT  X   MemberrZ  �r[  �r\  �r]  }r^  (hh]r_  �r`  Rra  hjW  uba�rb  Rrc  hh�jZ  j]  ubhhX   Functionrd  �re  �rf  �rg  }rh  (hh]ri  hhjd  h؇rj  �rk  �rl  }rm  (hh]rn  �ro  Rrp  hjg  uba�rq  Rrr  hh�h�jl  ubhhh�rs  �rt  �ru  }rv  (hh]rw  �rx  Rry  hh�ubhhh2�rz  �r{  �r|  }r}  (hh]r~  �r  Rr�  hh�ube�r�  Rr�  hh]h�h�j6  j9  h�h�h2j|  h�h�h�h�h�h�jd  jg  j  j  j'  j*  h:j  jT  jW  h�h�h�h�jL  jO  j  j  hBj"  hhj1  j  j  hju  ubhX   Literalr�  �r�  �r�  �r�  }r�  (hh]r�  (hj�  jT  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hj�  ubhj�  X   Charr�  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hj�  ubhj�  X   Dater�  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hj�  ubhj�  X   Scalarr�  �r�  �r�  �r�  }r�  (hh]r�  hj�  j�  X   Plainr�  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hj�  uba�r�  Rr�  hj�  j�  j�  ubhj�  X   Stringr�  �r�  �r�  �r�  }r�  (hh]r�  (hj�  j�  X   Interpolr�  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hj�  ubhj�  j�  X	   Delimeterr�  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hj�  ubhj�  j�  j�  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hj�  ubhj�  j�  j  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hj�  ubhj�  j�  X   Singler�  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hj�  ubhj�  j�  jT  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hj�  ubhj�  j�  X   Backtickr�  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hj�  ubhj�  j�  h`�r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hj�  ubhj�  j�  X   Regexr�  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hj�  ubhj�  j�  X   Momentr�  �r�  �r�  �r�  }r�  (hh]r�  �r   Rr  hj�  ubhj�  j�  X   Booleanr  �r  �r  �r  }r  (hh]r  �r  Rr	  hj�  ubhj�  j�  X	   Characterr
  �r  �r  �r  }r  (hh]r  �r  Rr  hj�  ubhj�  j�  X	   Delimiterr  �r  �r  �r  }r  (hh]r  �r  Rr  hj�  ubhj�  j�  X   Docr  �r  �r  �r  }r  (hh]r  �r   Rr!  hj�  ubhj�  j�  h�r"  �r#  �r$  }r%  (hh]r&  �r'  Rr(  hj�  ubhj�  j�  X   Affixr)  �r*  �r+  �r,  }r-  (hh]r.  �r/  Rr0  hj�  ubhj�  j�  X   Heredocr1  �r2  �r3  �r4  }r5  (hh]r6  �r7  Rr8  hj�  ubhj�  j�  X   Doubler9  �r:  �r;  �r<  }r=  (hh]r>  �r?  Rr@  hj�  ubhj�  j�  X   InterprA  �rB  �rC  �rD  }rE  (hh]rF  �rG  RrH  hj�  ubhj�  j�  X   AtomrI  �rJ  �rK  �rL  }rM  (hh]rN  �rO  RrP  hj�  ube�rQ  RrR  hj�  j)  j,  j�  j�  j�  j�  j  j  j  j  j9  j<  h`j�  j1  j4  j�  j�  jT  j�  j�  j�  j�  j�  j  j�  j
  j  j�  j�  jA  jD  j  j  j�  j�  jI  jL  hj$  ubhj�  X   NumberrS  �rT  �rU  �rV  }rW  (hh]rX  (hj�  jS  X   FloatrY  �rZ  �r[  �r\  }r]  (hh]r^  �r_  Rr`  hjV  ubhj�  jS  X   Decra  �rb  �rc  �rd  }re  (hh]rf  �rg  Rrh  hjV  ubhj�  jS  X   Radixri  �rj  �rk  �rl  }rm  (hh]rn  �ro  Rrp  hjV  ubhj�  jS  X   Octrq  �rr  �rs  �rt  }ru  (hh]rv  �rw  Rrx  hjV  ubhj�  jS  X   Binry  �rz  �r{  �r|  }r}  (hh]r~  �r  Rr�  hjV  ubhj�  jS  h�r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hjV  ubhj�  jS  X   Hexr�  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hjV  ubhj�  jS  X   Integerr�  �r�  �r�  �r�  }r�  (hh]r�  h(j�  jS  j�  X   Longr�  tr�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hj�  uba�r�  Rr�  hjV  j�  j�  ubhj�  jS  X   Decimalr�  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hjV  ube�r�  Rr�  hj�  jy  j|  jY  j\  j�  j�  j�  j�  jq  jt  ji  jl  h�j�  j�  j�  ja  jd  ube�r�  Rr�  hh]j�  j�  jS  jV  j�  j�  j�  j�  jT  j�  j�  j�  ubhX   Genericr�  �r�  �r�  �r�  }r�  (hh]r�  (hj�  X   Errorr�  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hj�  ubhj�  X
   Subheadingr�  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hj�  ubhj�  X	   Tracebackr�  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hj�  ubhj�  X   Outputr�  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hj�  ubhj�  X   Promptr�  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hj�  ubhj�  X   Deletedr�  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hj�  ubhj�  X   Insertedr�  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hj�  ubhj�  X   Headingr�  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hj�  ubhj�  X   Strongr�  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hj�  ubhj�  X   Emphr�  �r�  �r�  �r�  }r�  (hh]r�  �r   Rr  hj�  ube�r  Rr  hh]j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  ubhj�  �r  �r  �r  }r  (hh]r  �r	  Rr
  hh]ubhhjT  �r  �r  �r  }r  (hh]r  �r  Rr  hh]ubhX   Textr  �r  �r  �r  }r  (hh]r  (hj  X   Rootr  �r  �r  �r  }r  (hh]r  �r  Rr  hj  ubhj  j  �r   �r!  �r"  }r#  (hh]r$  �r%  Rr&  hj  ubhj  X   Ragr'  �r(  �r)  �r*  }r+  (hh]r,  �r-  Rr.  hj  ubhj  X
   Whitespacer/  �r0  �r1  �r2  }r3  (hh]r4  �r5  Rr6  hj  ubhj  X   Beerr7  �r8  �r9  �r:  }r;  (hh]r<  �r=  Rr>  hj  ubhj  X   Punctuationr?  �r@  �rA  �rB  }rC  (hh]rD  �rE  RrF  hj  ube�rG  RrH  hh]j/  j2  j  j"  j?  jB  j  j  j7  j:  j'  j*  ubhX   CommentrI  �rJ  �rK  �rL  }rM  (hh]rN  (hjI  X   PreprocrO  �rP  �rQ  �rR  }rS  (hh]rT  �rU  RrV  hjL  ubhjI  X   MultirW  �rX  �rY  �rZ  }r[  (hh]r\  �r]  Rr^  hjL  ubhjI  X   Hashbangr_  �r`  �ra  �rb  }rc  (hh]rd  �re  Rrf  hjL  ubhjI  j�  �rg  �rh  �ri  }rj  (hh]rk  �rl  Rrm  hjL  ubhjI  X
   SingleLinern  �ro  �rp  �rq  }rr  (hh]rs  �rt  Rru  hjL  ubhjI  j  �rv  �rw  �rx  }ry  (hh]rz  �r{  Rr|  hjL  ubhjI  X	   Directiver}  �r~  �r  �r�  }r�  (hh]r�  �r�  Rr�  hjL  ubhjI  X	   Multiliner�  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hjL  ubhjI  X
   Singleliner�  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hjL  ubhjI  X   PreprocFiler�  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hjL  ubhjI  X   Specialr�  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hjL  ube�r�  Rr�  hh]j_  jb  j�  j�  jO  jR  j�  j�  j�  ji  j�  j�  j}  j�  jn  jq  j  jx  jW  jZ  j�  j�  ubhj?  �r�  �r�  �r�  }r�  (hh]r�  hj?  X	   Indicatorr�  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hj�  uba�r�  Rr�  hh]j�  j�  ube�r�  Rr�  j  j  h`hcj�  j  jT  j  hhhh�j�  j�  j?  j�  hhhkjI  jL  j�  j�  X   Tokenr�  h]j�  j�  jS  jV  ubh2h5hJhMh:h=hBhEhRhUhhh*h-hhh"h%h
hubX   moduler�  �r�  j  X    r�  �r�  h�X   toplevelr�  �r�  j�  X   (r�  �r�  h�X   clockr�  �r�  j�  X   ,r�  �r�  h�X   resetr�  �r�  j�  X   )r�  �r�  j�  X   ;r�  �r�  j  X   
r�  �r�  j  j�  �r�  hX   inputr�  �r�  j  j�  �r�  h�X   clockr�  �r�  j�  j�  �r�  j  j�  �r�  j  j�  �r�  hX   inputr�  �r�  j  j�  �r�  h�X   resetr�  �r�  j�  j�  �r�  j  j�  �r�  j  X    
 r�  �r�  hX   regr�  �r�  j  j�  �r�  h�X   flop1r�  �r�  j�  j�  �r�  j  j�  �r�  j  j�  �r�  hX   regr�  �r�  j  j�  �r�  h�X   flop2r�  �r�  j�  j�  �r�  j  j�  �r�  j  X    
 r�  �r�  hX   alwaysr�  �r�  j  j�  �r�  j�  X   @r�  �r�  j  j�  �r�  j�  j�  �r�  hX   posedger�  �r�  j  j�  �r�  h�X   resetr�  �r�  j  j�  �r�  hX   orr�  �r�  j  j�  �r�  hX   posedger   �r  j  j�  �r  h�X   clockr  �r  j�  j�  �r  j  j�  �r  j  j�  �r  hX   ifr  �r	  j  j�  �r
  j�  j�  �r  h�X   resetr  �r  j�  j�  �r  j  j�  �r  j  X      r  �r  hX   beginr  �r  j  j�  �r  j  X        r  �r  h�X   flop1r  �r  j  j�  �r  hkX   <r  �r  hkX   =r  �r  j  j�  �r  j�  X   0r  �r   j�  j�  �r!  j  j�  �r"  j  X        r#  �r$  h�X   flop2r%  �r&  j  j�  �r'  hkj  �r(  hkj  �r)  j  j�  �r*  j�  X   1r+  �r,  j�  j�  �r-  j  j�  �r.  j  X      r/  �r0  hX   endr1  �r2  j  j�  �r3  j  j�  �r4  hX   elser5  �r6  j  j�  �r7  j  X      r8  �r9  hX   beginr:  �r;  j  j�  �r<  j  X        r=  �r>  h�X   flop1r?  �r@  j  j�  �rA  hkj  �rB  hkj  �rC  j  j�  �rD  h�X   flop2rE  �rF  j�  j�  �rG  j  j�  �rH  j  X        rI  �rJ  h�X   flop2rK  �rL  j  j�  �rM  hkj  �rN  hkj  �rO  j  j�  �rP  h�X   flop1rQ  �rR  j�  j�  �rS  j  j�  �rT  j  X      rU  �rV  hX   endrW  �rX  j  j�  �rY  hX	   endmodulerZ  �r[  j  j�  �r\  e.