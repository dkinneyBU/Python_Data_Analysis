�]q (cpygments.token
_TokenType
qX   Keywordq�q�q�q}q(X   subtypesqcbuiltins
set
q]q	(hhX   Wordq
�q�q�q}q(hh]q�qRqX   parentqhubhhh�q�q�q}q(hh]q�qRqhhubhhX   Typeq�q�q�q}q(hh]q�q Rq!hhubhhX   PreProcq"�q#�q$�q%}q&(hh]q'�q(Rq)hhubhhX   Controlq*�q+�q,�q-}q.(hh]q/�q0Rq1hhubhhX   Constantq2�q3�q4�q5}q6(hh]q7�q8Rq9hhubhhX	   Namespaceq:�q;�q<�q=}q>(hh]q?�q@RqAhhubhhX   PseudoqB�qC�qD�qE}qF(hh]qG�qHRqIhhubhhX   DeclarationqJ�qK�qL�qM}qN(hh]qO�qPRqQhhubhhX   ReservedqR�qS�qT�qU}qV(hh]qW�qXRqYhhube�qZRq[hh)�q\�q]}q^(hh]q_(hX   Escapeq`�qa�qb�qc}qd(hh]qe�qfRqghh]ubhX   Operatorqh�qi�qj�qk}ql(hh]qm(hhhX   DBSqn�qo�qp�qq}qr(hh]qs�qtRquhhkubhhhh
�qv�qw�qx}qy(hh]qz�q{Rq|hhkube�q}Rq~hh]h
hxhnhqubhX   Nameq�q��q��q�}q�(hh]q�(hhX   Tagq��q��q��q�}q�(hh]q��q�Rq�hh�ubhhX   Entityq��q��q��q�}q�(hh]q�hhh�hn�q��q��q�}q�(hh]q��q�Rq�hh�uba�q�Rq�hh�hnh�ubhhX	   Exceptionq��q��q��q�}q�(hh]q��q�Rq�hh�ubhhX	   Decoratorq��q��q��q�}q�(hh]q��q�Rq�hh�ubhhX   Classq��q��q��q�}q�(hh]q�(hhh�hn�q��q��q�}q�(hh]q��q�Rq�hh�ubhhh�X   Startq��q��q��q�}q�(hh]q��q�Rq�hh�ube�q�Rq�hh�h�h�hnh�ubhhX   VariableqÆqąqŁq�}q�(hh]q�(hhh�X	   Anonymousqɇqʅqˁq�}q�(hh]q΅q�Rq�hh�ubhhh�h��qхqҁq�}q�(hh]qՅq�Rq�hh�ubhhh�X   Magicq؇qمqځq�}q�(hh]q݅q�Rq�hh�ubhhh�X   Globalq��q�q�q�}q�(hh]q�q�Rq�hh�ubhhh�X   Instanceq�q�q�q�}q�(hh]q�q�Rq�hh�ube�q�Rq�hh�h�h�h�h�h�h�h�h�h�h�ubhhX	   Attributeq�q�q�q�}q�(hh]q�hhh�hÇq��q��q�}q�(hh]q��q�Rq�hh�uba�q�Rr   hh�h�h�ubhhh:�r  �r  �r  }r  (hh]r  �r  Rr  hh�ubhhX   Propertyr  �r	  �r
  �r  }r  (hh]r  �r  Rr  hh�ubhhX   Symbolr  �r  �r  �r  }r  (hh]r  �r  Rr  hh�ubhhX   Classesr  �r  �r  �r  }r  (hh]r  �r  Rr  hh�ubhhhB�r   �r!  �r"  }r#  (hh]r$  �r%  Rr&  hh�ubhhX   Labelr'  �r(  �r)  �r*  }r+  (hh]r,  �r-  Rr.  hh�ubhhhh�r/  �r0  �r1  }r2  (hh]r3  �r4  Rr5  hh�ubhhX   Builtinr6  �r7  �r8  �r9  }r:  (hh]r;  (hhj6  hB�r<  �r=  �r>  }r?  (hh]r@  �rA  RrB  hj9  ubhhj6  h�rC  �rD  �rE  }rF  (hh]rG  �rH  RrI  hj9  ube�rJ  RrK  hh�hBj>  hjE  ubhhX   FieldrL  �rM  �rN  �rO  }rP  (hh]rQ  �rR  RrS  hh�ubhhX   OtherrT  �rU  �rV  �rW  }rX  (hh]rY  hhjT  X   MemberrZ  �r[  �r\  �r]  }r^  (hh]r_  �r`  Rra  hjW  uba�rb  Rrc  hh�jZ  j]  ubhhX   Functionrd  �re  �rf  �rg  }rh  (hh]ri  hhjd  h؇rj  �rk  �rl  }rm  (hh]rn  �ro  Rrp  hjg  uba�rq  Rrr  hh�h�jl  ubhhh�rs  �rt  �ru  }rv  (hh]rw  �rx  Rry  hh�ubhhh2�rz  �r{  �r|  }r}  (hh]r~  �r  Rr�  hh�ube�r�  Rr�  hh]h�h�j6  j9  h�h�h2j|  h�h�h�h�h�h�jd  jg  j  j  j'  j*  h:j  jT  jW  h�h�h�h�jL  jO  j  j  hBj"  hhj1  j  j  hju  ubhX   Literalr�  �r�  �r�  �r�  }r�  (hh]r�  (hj�  jT  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hj�  ubhj�  X   Charr�  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hj�  ubhj�  X   Dater�  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hj�  ubhj�  X   Scalarr�  �r�  �r�  �r�  }r�  (hh]r�  hj�  j�  X   Plainr�  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hj�  uba�r�  Rr�  hj�  j�  j�  ubhj�  X   Stringr�  �r�  �r�  �r�  }r�  (hh]r�  (hj�  j�  X   Interpolr�  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hj�  ubhj�  j�  X	   Delimeterr�  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hj�  ubhj�  j�  j�  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hj�  ubhj�  j�  j  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hj�  ubhj�  j�  X   Singler�  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hj�  ubhj�  j�  jT  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hj�  ubhj�  j�  X   Backtickr�  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hj�  ubhj�  j�  h`�r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hj�  ubhj�  j�  X   Regexr�  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hj�  ubhj�  j�  X   Momentr�  �r�  �r�  �r�  }r�  (hh]r�  �r   Rr  hj�  ubhj�  j�  X   Booleanr  �r  �r  �r  }r  (hh]r  �r  Rr	  hj�  ubhj�  j�  X	   Characterr
  �r  �r  �r  }r  (hh]r  �r  Rr  hj�  ubhj�  j�  X	   Delimiterr  �r  �r  �r  }r  (hh]r  �r  Rr  hj�  ubhj�  j�  X   Docr  �r  �r  �r  }r  (hh]r  �r   Rr!  hj�  ubhj�  j�  h�r"  �r#  �r$  }r%  (hh]r&  �r'  Rr(  hj�  ubhj�  j�  X   Affixr)  �r*  �r+  �r,  }r-  (hh]r.  �r/  Rr0  hj�  ubhj�  j�  X   Heredocr1  �r2  �r3  �r4  }r5  (hh]r6  �r7  Rr8  hj�  ubhj�  j�  X   Doubler9  �r:  �r;  �r<  }r=  (hh]r>  �r?  Rr@  hj�  ubhj�  j�  X   InterprA  �rB  �rC  �rD  }rE  (hh]rF  �rG  RrH  hj�  ubhj�  j�  X   AtomrI  �rJ  �rK  �rL  }rM  (hh]rN  �rO  RrP  hj�  ube�rQ  RrR  hj�  j)  j,  j�  j�  j�  j�  j  j  j  j  j9  j<  h`j�  j1  j4  j�  j�  jT  j�  j�  j�  j�  j�  j  j�  j
  j  j�  j�  jA  jD  j  j  j�  j�  jI  jL  hj$  ubhj�  X   NumberrS  �rT  �rU  �rV  }rW  (hh]rX  (hj�  jS  X   FloatrY  �rZ  �r[  �r\  }r]  (hh]r^  �r_  Rr`  hjV  ubhj�  jS  X   Decra  �rb  �rc  �rd  }re  (hh]rf  �rg  Rrh  hjV  ubhj�  jS  X   Radixri  �rj  �rk  �rl  }rm  (hh]rn  �ro  Rrp  hjV  ubhj�  jS  X   Octrq  �rr  �rs  �rt  }ru  (hh]rv  �rw  Rrx  hjV  ubhj�  jS  X   Binry  �rz  �r{  �r|  }r}  (hh]r~  �r  Rr�  hjV  ubhj�  jS  h�r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hjV  ubhj�  jS  X   Hexr�  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hjV  ubhj�  jS  X   Integerr�  �r�  �r�  �r�  }r�  (hh]r�  h(j�  jS  j�  X   Longr�  tr�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hj�  uba�r�  Rr�  hjV  j�  j�  ubhj�  jS  X   Decimalr�  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hjV  ube�r�  Rr�  hj�  jy  j|  jY  j\  j�  j�  j�  j�  jq  jt  ji  jl  h�j�  j�  j�  ja  jd  ube�r�  Rr�  hh]j�  j�  jS  jV  j�  j�  j�  j�  jT  j�  j�  j�  ubhX   Genericr�  �r�  �r�  �r�  }r�  (hh]r�  (hj�  X   Errorr�  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hj�  ubhj�  X
   Subheadingr�  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hj�  ubhj�  X	   Tracebackr�  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hj�  ubhj�  X   Outputr�  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hj�  ubhj�  X   Promptr�  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hj�  ubhj�  X   Deletedr�  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hj�  ubhj�  X   Insertedr�  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hj�  ubhj�  X   Headingr�  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hj�  ubhj�  X   Strongr�  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hj�  ubhj�  X   Emphr�  �r�  �r�  �r�  }r�  (hh]r�  �r   Rr  hj�  ube�r  Rr  hh]j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  ubhj�  �r  �r  �r  }r  (hh]r  �r	  Rr
  hh]ubhhjT  �r  �r  �r  }r  (hh]r  �r  Rr  hh]ubhX   Textr  �r  �r  �r  }r  (hh]r  (hj  X   Rootr  �r  �r  �r  }r  (hh]r  �r  Rr  hj  ubhj  j  �r   �r!  �r"  }r#  (hh]r$  �r%  Rr&  hj  ubhj  X   Ragr'  �r(  �r)  �r*  }r+  (hh]r,  �r-  Rr.  hj  ubhj  X
   Whitespacer/  �r0  �r1  �r2  }r3  (hh]r4  �r5  Rr6  hj  ubhj  X   Beerr7  �r8  �r9  �r:  }r;  (hh]r<  �r=  Rr>  hj  ubhj  X   Punctuationr?  �r@  �rA  �rB  }rC  (hh]rD  �rE  RrF  hj  ube�rG  RrH  hh]j/  j2  j  j"  j?  jB  j  j  j7  j:  j'  j*  ubhX   CommentrI  �rJ  �rK  �rL  }rM  (hh]rN  (hjI  X   PreprocrO  �rP  �rQ  �rR  }rS  (hh]rT  �rU  RrV  hjL  ubhjI  X   MultirW  �rX  �rY  �rZ  }r[  (hh]r\  �r]  Rr^  hjL  ubhjI  X   Hashbangr_  �r`  �ra  �rb  }rc  (hh]rd  �re  Rrf  hjL  ubhjI  j�  �rg  �rh  �ri  }rj  (hh]rk  �rl  Rrm  hjL  ubhjI  X
   SingleLinern  �ro  �rp  �rq  }rr  (hh]rs  �rt  Rru  hjL  ubhjI  j  �rv  �rw  �rx  }ry  (hh]rz  �r{  Rr|  hjL  ubhjI  X	   Directiver}  �r~  �r  �r�  }r�  (hh]r�  �r�  Rr�  hjL  ubhjI  X	   Multiliner�  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hjL  ubhjI  X
   Singleliner�  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hjL  ubhjI  X   PreprocFiler�  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hjL  ubhjI  X   Specialr�  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hjL  ube�r�  Rr�  hh]j_  jb  j�  j�  jO  jR  j�  j�  j�  ji  j�  j�  j}  j�  jn  jq  j  jx  jW  jZ  j�  j�  ubhj?  �r�  �r�  �r�  }r�  (hh]r�  hj?  X	   Indicatorr�  �r�  �r�  �r�  }r�  (hh]r�  �r�  Rr�  hj�  uba�r�  Rr�  hh]j�  j�  ube�r�  Rr�  j  j  h`hcj�  j  jT  j  hhhh�j�  j�  j?  j�  hhhkjI  jL  j�  j�  X   Tokenr�  h]j�  j�  jS  jV  ubh2h5hJhMh:h=hBhEhRhUhhh*h-hhh"h%h
hubX   libraryr�  �r�  j  X    r�  �r�  j  X   ieeer�  �r�  j�  X   ;r�  �r�  j  X   
r�  �r�  hX   user�  �r�  j  j�  �r�  j  X   ieee.std_logic_unsigned.r�  �r�  hX   allr�  �r�  j�  j�  �r�  j  j�  �r�  hX   user�  �r�  j  j�  �r�  j  X   ieee.std_logic_1164.r�  �r�  hX   allr�  �r�  j�  j�  �r�  j  X      
r�  �r�  hX   user�  �r�  j  j�  �r�  j  X   ieee.numeric_std.r�  �r�  hX   allr�  �r�  j�  j�  �r�  j  j�  �r�  j  j�  �r�  j  j�  �r�  hX   entityr�  �r�  j  j�  �r�  h�X   top_testbenchr�  �r�  j  j�  �r�  hX   isr�  �r�  j  j�  �r�  ji  X   --testr�  �r�  j  j�  �r�  j  X   	r�  �r�  hX   genericr�  �r�  j  j�  �r�  j�  X   (r�  �r�  j  j�  �r�  ji  X   -- testr�  �r�  j  j�  �r�  j  X   	    r�  �r�  h�X   nr�  �r�  j  j�  �r�  hkX   :r�  �r�  j  j�  �r�  hX   integerr   �r  j  j�  �r  hkj�  �r  hkX   =r  �r  j  j�  �r  j�  X   8r  �r  j  j�  �r	  ji  X   -- testr
  �r  j  j�  �r  j  j�  �r  j�  X   )r  �r  j�  j�  �r  j  j�  �r  ji  X   -- testr  �r  j  j�  �r  hX   endr  �r  j  j�  �r  h�X   top_testbenchr  �r  j�  j�  �r  j  j�  �r  ji  X   -- testr  �r  j  j�  �r  j  j�  �r  j  j�  �r   hX   architecturer!  �r"  j  j�  �r#  h�X   top_testbench_archr$  �r%  j  j�  �r&  hX   ofr'  �r(  j  j�  �r)  h�X   top_testbenchr*  �r+  j  j�  �r,  hX   isr-  �r.  j  X     

    r/  �r0  hX	   componentr1  �r2  j  j�  �r3  h�X   topr4  �r5  j  j�  �r6  hX   isr7  �r8  j  j�  �r9  j  X           r:  �r;  hX   genericr<  �r=  j  j�  �r>  j�  j�  �r?  j  j�  �r@  j  X               rA  �rB  h�j�  �rC  j  j�  �rD  hkj�  �rE  j  j�  �rF  hX   integerrG  �rH  j  j�  �rI  j  X           rJ  �rK  j�  j  �rL  j  X      rM  �rN  j�  j�  �rO  j  j�  �rP  j  X           rQ  �rR  hX   portrS  �rT  j  j�  �rU  j�  j�  �rV  j  j�  �rW  j  X               rX  �rY  h�X   clkrZ  �r[  j  j�  �r\  hkj�  �r]  j  j�  �r^  hX   inr_  �r`  j  j�  �ra  hX	   std_logicrb  �rc  j�  j�  �rd  j  j�  �re  j  X               rf  �rg  h�X   rstrh  �ri  j  j�  �rj  hkj�  �rk  j  j�  �rl  hX   inrm  �rn  j  j�  �ro  hX	   std_logicrp  �rq  j�  j�  �rr  j  j�  �rs  j  X               rt  �ru  h�X   d1rv  �rw  j  j�  �rx  hkj�  �ry  j  j�  �rz  hX   inr{  �r|  j  j�  �r}  hX   std_logic_vectorr~  �r  j  j�  �r�  j�  j�  �r�  h�j�  �r�  hkX   -r�  �r�  j�  X   1r�  �r�  j  j�  �r�  hX   downtor�  �r�  j  j�  �r�  j�  X   0r�  �r�  j�  j  �r�  j�  j�  �r�  j  j�  �r�  j  X               r�  �r�  h�X   d2r�  �r�  j  j�  �r�  hkj�  �r�  j  j�  �r�  hX   inr�  �r�  j  j�  �r�  hX   std_logic_vectorr�  �r�  j  j�  �r�  j�  j�  �r�  h�j�  �r�  hkj�  �r�  j�  j�  �r�  j  j�  �r�  hX   downtor�  �r�  j  j�  �r�  j�  j�  �r�  j�  j  �r�  j�  j�  �r�  j  j�  �r�  j  X               r�  �r�  h�X	   operationr�  �r�  j  j�  �r�  hkj�  �r�  j  j�  �r�  hX   inr�  �r�  j  j�  �r�  hX	   std_logicr�  �r�  j�  j�  �r�  j  j�  �r�  j  X               r�  �r�  h�X   resultr�  �r�  j  j�  �r�  hkj�  �r�  j  j�  �r�  hX   outr�  �r�  j  j�  �r�  hX   std_logic_vectorr�  �r�  j  j�  �r�  j�  j�  �r�  j�  X   2r�  �r�  hkX   *r�  �r�  h�j�  �r�  hkj�  �r�  j�  j�  �r�  j  j�  �r�  hX   downtor�  �r�  j  j�  �r�  j�  j�  �r�  j�  j  �r�  j  j�  �r�  j  X           r�  �r�  j�  j  �r�  j�  j�  �r�  j  j�  �r�  j  X       r�  �r�  hX   endr�  �r�  j  j�  �r�  hX	   componentr�  �r�  j�  j�  �r�  j  j�  �r�  j  j�  �r�  j  X       r�  �r�  hX   signalr�  �r�  j  j�  �r�  h�X   clkr�  �r�  j  j�  �r�  hkj�  �r�  j  j�  �r�  hX	   std_logicr�  �r�  j�  j�  �r�  j  j�  �r�  j  X       r�  �r�  hX   signalr�  �r�  j  j�  �r�  h�X   rstr�  �r�  j  j�  �r�  hkj�  �r�  j  j�  �r�  hX	   std_logicr�  �r�  j�  j�  �r�  j  j�  �r�  j  j�  �r�  hX   signalr�  �r   j  j�  �r  h�X	   operationr  �r  j  j�  �r  hkj�  �r  j  j�  �r  hX	   std_logicr  �r  j�  j�  �r	  j  j�  �r
  j  X       r  �r  hX   signalr  �r  j  j�  �r  h�X   d1r  �r  j  j�  �r  hkj�  �r  j  j�  �r  hX   std_logic_vectorr  �r  j  j�  �r  j�  j�  �r  h�j�  �r  hkj�  �r  j�  j�  �r  j  j�  �r  hX   downtor  �r  j  j�  �r  j�  j�  �r   j�  j  �r!  j�  j�  �r"  j  j�  �r#  j  X       r$  �r%  hX   signalr&  �r'  j  j�  �r(  h�X   d2r)  �r*  j  j�  �r+  hkj�  �r,  j  j�  �r-  hX   std_logic_vectorr.  �r/  j  j�  �r0  j�  j�  �r1  h�j�  �r2  hkj�  �r3  j�  j�  �r4  j  j�  �r5  hX   downtor6  �r7  j  j�  �r8  j�  j�  �r9  j�  j  �r:  j�  j�  �r;  j  j�  �r<  j  X       r=  �r>  hX   signalr?  �r@  j  j�  �rA  h�X   resultrB  �rC  j  j�  �rD  hkj�  �rE  j  j�  �rF  hX   std_logic_vectorrG  �rH  j  j�  �rI  j�  j�  �rJ  j�  j�  �rK  hkj�  �rL  h�j�  �rM  hkj�  �rN  j�  j�  �rO  j  j�  �rP  hX   downtorQ  �rR  j  j�  �rS  j�  j�  �rT  j�  j  �rU  j�  j�  �rV  j  j�  �rW  j  X	       
    rX  �rY  hX   typerZ  �r[  j  j�  �r\  h�X	   test_typer]  �r^  j  j�  �r_  hX   isr`  �ra  j  j�  �rb  j�  j�  �rc  j  j�  �rd  h�X   a1re  �rf  j�  X   ,rg  �rh  j  j�  �ri  h�X   a2rj  �rk  j�  jg  �rl  j  j�  �rm  h�X   a3rn  �ro  j�  jg  �rp  j  j�  �rq  h�X   a4rr  �rs  j�  jg  �rt  j  j�  �ru  h�X   a5rv  �rw  j�  jg  �rx  j  j�  �ry  h�X   a6rz  �r{  j�  jg  �r|  j  j�  �r}  h�X   a7r~  �r  j�  jg  �r�  j  j�  �r�  h�X   a8r�  �r�  j�  jg  �r�  j  j�  �r�  h�X   a9r�  �r�  j�  jg  �r�  j  j�  �r�  h�X   a10r�  �r�  j�  j  �r�  j�  j�  �r�  j  j�  �r�  j  X       r�  �r�  hX	   attributer�  �r�  j  j�  �r�  h�X   enum_encodingr�  �r�  j  j�  �r�  hX   ofr�  �r�  j  j�  �r�  h�X   my_stater�  �r�  j  j�  �r�  hkj�  �r�  j  j�  �r�  hX   typer�  �r�  j  j�  �r�  hX   isr�  �r�  j  j�  �r�  j�  X   "001 010 011 100 111"r�  �r�  j�  j�  �r�  j  j�  �r�  hX   beginr�  �r�  j  j�  �r�  j  j�  �r�  j  X       r�  �r�  h�X   TESTUNITr�  �r�  j  j�  �r�  hkj�  �r�  j  j�  �r�  h�X   topr�  �r�  j  j�  �r�  hX   genericr�  �r�  j  j�  �r�  hX   mapr�  �r�  j  j�  �r�  j�  j�  �r�  h�j�  �r�  j  j�  �r�  hkj  �r�  hkX   >r�  �r�  j  j�  �r�  h�j�  �r�  j�  j  �r�  j  j�  �r�  j  X                      r�  �r�  hX   portr�  �r�  j  j�  �r�  hX   mapr�  �r�  j  j�  �r�  j�  j�  �r�  h�X   clkr�  �r�  j  j�  �r�  hkj  �r�  hkj�  �r�  j  j�  �r�  h�X   clkr�  �r�  j�  jg  �r�  j  j�  �r�  j  X                                r�  �r�  h�X   rstr�  �r�  j  j�  �r�  hkj  �r�  hkj�  �r�  j  j�  �r�  h�X   rstr�  �r�  j�  jg  �r�  j  j�  �r�  j  X                                r�  �r�  h�X   d1r�  �r�  j  X     r�  �r�  hkj  �r�  hkj�  �r�  j  j�  �r�  h�X   d1r�  �r�  j�  jg  �r�  j  j�  �r�  j  X                                r�  �r�  h�X   d2r�  �r�  j  X     r�  �r�  hkj  �r�  hkj�  �r�  j  j�  �r�  h�X   d2r�  �r�  j�  jg  �r�  j  j�  �r�  j  X                                r   �r  h�X	   operationr  �r  j  j�  �r  hkj  �r  hkj�  �r  j  j�  �r  h�X	   operationr  �r	  j�  jg  �r
  j  j�  �r  j  X                                r  �r  h�X   resultr  �r  j  j�  �r  hkj  �r  hkj�  �r  j  j�  �r  h�X   resultr  �r  j�  j  �r  j�  j�  �r  j  j�  �r  j  j�  �r  j  X       r  �r  h�X   clock_processr  �r  j  j�  �r  hkj�  �r  j  j�  �r   hX   processr!  �r"  j  j�  �r#  j  X       r$  �r%  hX   beginr&  �r'  j  j�  �r(  j  X           r)  �r*  h�X   clkr+  �r,  j  j�  �r-  hkX   <r.  �r/  hkj  �r0  j  j�  �r1  j�  X   '0'r2  �r3  j�  j�  �r4  j  j�  �r5  j  X           r6  �r7  hX   waitr8  �r9  j  j�  �r:  hX   forr;  �r<  j  j�  �r=  j�  X   5r>  �r?  j  j�  �r@  h�X   nsrA  �rB  j�  j�  �rC  j  j�  �rD  j  X           rE  �rF  h�X   clkrG  �rH  j  j�  �rI  hkj.  �rJ  hkj  �rK  j  j�  �rL  j�  X   '1'rM  �rN  j�  j�  �rO  j  j�  �rP  j  X           rQ  �rR  hX   waitrS  �rT  j  j�  �rU  hX   forrV  �rW  j  j�  �rX  j�  j>  �rY  j  j�  �rZ  h�X   nsr[  �r\  j�  j�  �r]  j  j�  �r^  j  X       r_  �r`  hX   endra  �rb  j  j�  �rc  hX   processrd  �re  j�  j�  �rf  j  j�  �rg  j  j�  �rh  j  X       ri  �rj  h�X   data_processrk  �rl  j  j�  �rm  hkj�  �rn  j  j�  �ro  hX   processrp  �rq  j  j�  �rr  j  X       rs  �rt  hX   beginru  �rv  j  X          
		
		rw  �rx  ji  X   -- test case #1	ry  �rz  j  j�  �r{  j  X   	   	r|  �r}  h�X	   operationr~  �r  j  j�  �r�  hkj.  �r�  hkj  �r�  j  j�  �r�  j�  X   '0'r�  �r�  j�  j�  �r�  j  j�  �r�  j  X   		
        r�  �r�  h�X   rstr�  �r�  j  j�  �r�  hkj.  �r�  hkj  �r�  j  j�  �r�  j�  X   '1'r�  �r�  j�  j�  �r�  j  j�  �r�  j  X           r�  �r�  hX   waitr�  �r�  j  j�  �r�  hX   forr�  �r�  j  j�  �r�  j�  j>  �r�  j  j�  �r�  h�X   nsr�  �r�  j�  j�  �r�  j  j�  �r�  j  X           r�  �r�  h�X   rstr�  �r�  j  j�  �r�  hkj.  �r�  hkj  �r�  j  j�  �r�  j�  X   '0'r�  �r�  j�  j�  �r�  j  j�  �r�  j  X           r�  �r�  hX   waitr�  �r�  j  j�  �r�  hX   forr�  �r�  j  j�  �r�  j�  j>  �r�  j  j�  �r�  h�X   nsr�  �r�  j�  j�  �r�  j  j�  �r�  j  X   		
		r�  �r�  h�X   d1r�  �r�  j  j�  �r�  hkj.  �r�  hkj  �r�  j  j�  �r�  hX   std_logic_vectorr�  �r�  j�  j�  �r�  h�X   to_unsignedr�  �r�  j�  j�  �r�  j�  X   60r�  �r�  j�  jg  �r�  j  j�  �r�  h�X   d1r�  �r�  h�X   'lengthr�  �r�  j�  j  �r�  j�  j  �r�  j�  j�  �r�  j  j�  �r�  j  X   		r�  �r�  h�X   d2r�  �r�  j  j�  �r�  hkj.  �r�  hkj  �r�  j  j�  �r�  hX   std_logic_vectorr�  �r�  j�  j�  �r�  h�X   to_unsignedr�  �r�  j�  j�  �r�  j�  X   12r�  �r�  j�  jg  �r�  j  j�  �r�  h�X   d2r�  �r�  h�X   'lengthr�  �r�  j�  j  �r�  j�  j  �r�  j�  j�  �r�  j  j�  �r�  j  X   		r�  �r�  hX   waitr�  �r�  j  j�  �r�  hX   forr�  �r�  j  j�  �r�  j�  X   360r�  �r�  j  j�  �r�  h�X   nsr�  �r�  j�  j�  �r�  j  j�  �r�  j  X   		
		r�  �r   hX   assertr  �r  j  j�  �r  j�  j�  �r  h�X   resultr  �r  j  j�  �r  hkj  �r  j  j�  �r	  hX   std_logic_vectorr
  �r  j�  j�  �r  h�X   to_unsignedr  �r  j�  j�  �r  j�  X   720r  �r  j�  jg  �r  j  j�  �r  h�X   resultr  �r  h�X   'lengthr  �r  j�  j  �r  j�  j  �r  j�  j  �r  j  j�  �r  j  X   			r  �r  h�X   reportr  �r  j  j�  �r   j�  X   "Test case #1 failed"r!  �r"  j  j�  �r#  hX   severityr$  �r%  j  j�  �r&  h�X   errorr'  �r(  j�  j�  �r)  j  X    
            
		r*  �r+  ji  X   -- test case #2	r,  �r-  j  j�  �r.  j  X   	   	r/  �r0  h�X	   operationr1  �r2  j  j�  �r3  hkj.  �r4  hkj  �r5  j  j�  �r6  j�  X   '0'r7  �r8  j�  j�  �r9  j  j�  �r:  j  X   		
        r;  �r<  h�X   rstr=  �r>  j  j�  �r?  hkj.  �r@  hkj  �rA  j  j�  �rB  j�  X   '1'rC  �rD  j�  j�  �rE  j  j�  �rF  j  X           rG  �rH  hX   waitrI  �rJ  j  j�  �rK  hX   forrL  �rM  j  j�  �rN  j�  j>  �rO  j  j�  �rP  h�X   nsrQ  �rR  j�  j�  �rS  j  j�  �rT  j  X           rU  �rV  h�X   rstrW  �rX  j  j�  �rY  hkj.  �rZ  hkj  �r[  j  j�  �r\  j�  X   '0'r]  �r^  j�  j�  �r_  j  j�  �r`  j  X           ra  �rb  hX   waitrc  �rd  j  j�  �re  hX   forrf  �rg  j  j�  �rh  j�  j>  �ri  j  j�  �rj  h�X   nsrk  �rl  j�  j�  �rm  j  j�  �rn  j  X   		
		ro  �rp  h�X   d1rq  �rr  j  j�  �rs  hkj.  �rt  hkj  �ru  j  j�  �rv  hX   std_logic_vectorrw  �rx  j�  j�  �ry  h�X   to_unsignedrz  �r{  j�  j�  �r|  j�  X   55r}  �r~  j�  jg  �r  j  j�  �r�  h�X   d1r�  �r�  h�X   'lengthr�  �r�  j�  j  �r�  j�  j  �r�  j�  j�  �r�  j  j�  �r�  j  X   		r�  �r�  h�X   d2r�  �r�  j  j�  �r�  hkj.  �r�  hkj  �r�  j  j�  �r�  hX   std_logic_vectorr�  �r�  j�  j�  �r�  h�X   to_unsignedr�  �r�  j�  j�  �r�  j�  j�  �r�  j�  jg  �r�  j  j�  �r�  h�X   d2r�  �r�  h�X   'lengthr�  �r�  j�  j  �r�  j�  j  �r�  j�  j�  �r�  j  j�  �r�  j  X   		r�  �r�  hX   waitr�  �r�  j  j�  �r�  hX   forr�  �r�  j  j�  �r�  j�  X   360r�  �r�  j  j�  �r�  h�X   nsr�  �r�  j�  j�  �r�  j  j�  �r�  j  X   		
		r�  �r�  hX   assertr�  �r�  j  j�  �r�  j�  j�  �r�  h�X   resultr�  �r�  j  j�  �r�  hkj  �r�  j  j�  �r�  hX   std_logic_vectorr�  �r�  j�  j�  �r�  h�X   to_unsignedr�  �r�  j�  j�  �r�  j�  X   55r�  �r�  j�  jg  �r�  j  j�  �r�  h�X   resultr�  �r�  h�X   'lengthr�  �r�  j�  j  �r�  j�  j  �r�  j�  j  �r�  j  j�  �r�  j  X   			r�  �r�  h�X   reportr�  �r�  j  j�  �r�  j�  X   "Test case #2 failed"r�  �r�  j  j�  �r�  hX   severityr�  �r�  j  j�  �r�  h�X   errorr�  �r�  j�  j�  �r�  j  j�  �r�  j  X               
        r�  �r�  ji  X   -- etc r�  �r�  j  j�  �r�  j  X               
    r�  �r�  hX   endr�  �r�  j  j�  �r�  hX   processr�  �r�  j�  j�  �r�  j  j�  �r�  j  j�  �r�  hX   endr�  �r�  j  j�  �r�  h�X   top_testbench_archr�  �r�  j�  j�  �r�  j  j�  �r�  j  j�  �r�  j  j�  �r�  hX   configurationr�  �r�  j  j�  �r�  h�X   testbench_for_topr�  �r�  j  j�  �r�  hX   ofr�  �r�  j  j�  �r�  h�X   top_testbenchr�  �r�  j  j�  �r   hX   isr  �r  j  j�  �r  j  j�  �r  hX   forr  �r  j  j�  �r  h�X   top_testbench_archr  �r	  j  j�  �r
  j  X   		r  �r  hX   forr  �r  j  j�  �r  h�X   TESTUNITr  �r  j  j�  �r  hkj�  �r  j  j�  �r  h�X   topr  �r  j  j�  �r  j  X   			r  �r  hX   user  �r  j  j�  �r  hX   entityr  �r  j  j�  �r  j  X   workr   �r!  j�  X   .r"  �r#  h�X   topr$  �r%  j�  j�  �r&  h�X   top_archr'  �r(  j�  j  �r)  j�  j�  �r*  j  j�  �r+  j  X   		r,  �r-  hX   endr.  �r/  j  j�  �r0  hX   forr1  �r2  j�  j�  �r3  j  j�  �r4  j  j�  �r5  hX   endr6  �r7  j  j�  �r8  hX   forr9  �r:  j�  j�  �r;  j  j�  �r<  hX   endr=  �r>  j  j�  �r?  h�X   testbench_for_topr@  �rA  j�  j�  �rB  j  j�  �rC  j  j�  �rD  j  j�  �rE  hX   functionrF  �rG  j  j�  �rH  h�X   comparerI  �rJ  j�  j�  �rK  h�X   ArL  �rM  hkj�  �rN  j  j�  �rO  hX	   std_logicrP  �rQ  j�  jg  �rR  j  j�  �rS  h�X   BrT  �rU  hkj�  �rV  j  j�  �rW  hX	   std_LogicrX  �rY  j�  j  �rZ  j  j�  �r[  hX   returnr\  �r]  j  j�  �r^  hX	   std_logicr_  �r`  j  j�  �ra  hX   isrb  �rc  j  j�  �rd  j  X       re  �rf  hX   constantrg  �rh  j  j�  �ri  h�X   pirj  �rk  j  j�  �rl  hkj�  �rm  j  j�  �rn  h�X   realro  �rp  j  j�  �rq  hkj�  �rr  hkj  �rs  j  j�  �rt  j�  X   3ru  �rv  j�  j"  �rw  j�  X   14159rx  �ry  j�  j�  �rz  j  j�  �r{  j  X       r|  �r}  hX   constantr~  �r  j  j�  �r�  h�X   half_pir�  �r�  j  j�  �r�  hkj�  �r�  j  j�  �r�  h�X   realr�  �r�  j  j�  �r�  hkj�  �r�  hkj  �r�  j  j�  �r�  h�X   pir�  �r�  j  j�  �r�  hkX   /r�  �r�  j  j�  �r�  j�  j�  �r�  j�  j"  �r�  j�  j�  �r�  j�  j�  �r�  j  j�  �r�  j  X       r�  �r�  hX   constantr�  �r�  j  j�  �r�  h�X
   cycle_timer�  �r�  j  j�  �r�  hkj�  �r�  j  j�  �r�  hX   timer�  �r�  j  j�  �r�  hkj�  �r�  hkj  �r�  j  j�  �r�  j�  j�  �r�  j  j�  �r�  h�X   nsr�  �r�  j�  j�  �r�  j  j�  �r�  j  X       r�  �r�  hX   constantr�  �r�  j  j�  �r�  h�X   Nr�  �r�  j�  jg  �r�  j  j�  �r�  h�X   N5r�  �r�  j  j�  �r�  hkj�  �r�  j  j�  �r�  hX   integerr�  �r�  j  j�  �r�  hkj�  �r�  hkj  �r�  j  j�  �r�  j�  j>  �r�  j�  j�  �r�  j  j�  �r�  hX   beginr�  �r�  j  j�  �r�  j  X       r�  �r�  hX   ifr�  �r�  j  j�  �r�  j�  j�  �r�  h�jL  �r�  j  j�  �r�  hkj  �r�  j  j�  �r�  j�  X   '0'r�  �r�  j  j�  �r�  hX   andr�  �r�  j  j�  �r�  h�jT  �r�  j  j�  �r�  hkj  �r�  j  j�  �r�  j�  X   '1'r�  �r�  j�  j  �r�  j  j�  �r�  hX   thenr�  �r�  j  j�  �r�  j  X           r�  �r�  hX   returnr�  �r�  j  j�  �r�  h�jT  �r�  j�  j�  �r�  j  j�  �r�  j  X       r�  �r�  hX   elser�  �r�  j  j�  �r�  j  X           r�  �r�  hX   returnr�  �r�  j  j�  �r�  h�jL  �r�  j�  j�  �r�  j  j�  �r�  j  X       r�  �r�  hX   endr�  �r�  j  j�  �r�  hX   ifr�  �r�  j  j�  �r�  j�  j�  �r�  j  j�  �r 	  hX   endr	  �r	  j  j�  �r	  h�X   comparer	  �r	  j�  j�  �r	  j  j�  �r	  j  j�  �r	  j  j�  �r		  hX	   procedurer
	  �r	  j  j�  �r	  h�X   printr	  �r	  j�  j�  �r	  h�X   Pr	  �r	  j  j�  �r	  hkj�  �r	  j  j�  �r	  hX   std_logic_vectorr	  �r	  j�  j�  �r	  j�  X   7r	  �r	  j  j�  �r	  hX   downtor	  �r	  j  j�  �r	  j�  j�  �r	  j�  j  �r	  e(j�  j�  �r 	  j  j�  �r!	  j  X                   r"	  �r#	  h�X   Ur$	  �r%	  j  j�  �r&	  hkj�  �r'	  j  j�  �r(	  hX   std_logic_vectorr)	  �r*	  j�  j�  �r+	  j�  ju  �r,	  j  j�  �r-	  hX   downtor.	  �r/	  j  j�  �r0	  j�  j�  �r1	  j�  j  �r2	  j�  j  �r3	  j  j�  �r4	  hX   isr5	  �r6	  j  j�  �r7	  j  X       r8	  �r9	  hX   variabler:	  �r;	  j  j�  �r<	  h�X   my_liner=	  �r>	  j  j�  �r?	  hkj�  �r@	  j  j�  �rA	  h�X   linerB	  �rC	  j�  j�  �rD	  j  j�  �rE	  j  X       rF	  �rG	  hX   aliasrH	  �rI	  j  j�  �rJ	  h�X   swriterK	  �rL	  j  j�  �rM	  hX   isrN	  �rO	  j  j�  �rP	  h�X   writerQ	  �rR	  j  j�  �rS	  j�  X   [rT	  �rU	  h�X   linerV	  �rW	  j�  jg  �rX	  j  j�  �rY	  hX   stringrZ	  �r[	  j�  jg  �r\	  j  j�  �r]	  h�X   sider^	  �r_	  j�  jg  �r`	  j  j�  �ra	  h�X   widthrb	  �rc	  j�  X   ]rd	  �re	  j  j�  �rf	  j�  j�  �rg	  j  j�  �rh	  hX   beginri	  �rj	  j  j�  �rk	  j  X       rl	  �rm	  h�X   swritern	  �ro	  j�  j�  �rp	  h�X   my_linerq	  �rr	  j�  jg  �rs	  j  j�  �rt	  j�  X   "sqrt( "ru	  �rv	  j�  j  �rw	  j�  j�  �rx	  j  j�  �ry	  j  X       rz	  �r{	  h�X   writer|	  �r}	  j�  j�  �r~	  h�X   my_liner	  �r�	  j�  jg  �r�	  j  j�  �r�	  h�j	  �r�	  j�  j  �r�	  j�  j�  �r�	  j  j�  �r�	  j  X       r�	  �r�	  h�X   swriter�	  �r�	  j�  j�  �r�	  h�X   my_liner�	  �r�	  j�  jg  �r�	  j  j�  �r�	  j�  X   " )= "r�	  �r�	  j�  j  �r�	  j�  j�  �r�	  j  j�  �r�	  j  X       r�	  �r�	  h�X   writer�	  �r�	  j�  j�  �r�	  h�X   my_liner�	  �r�	  j�  jg  �r�	  j  j�  �r�	  h�j$	  �r�	  j�  j  �r�	  j�  j�  �r�	  j  j�  �r�	  j  X       r�	  �r�	  h�X	   writeliner�	  �r�	  j�  j�  �r�	  h�X   outputr�	  �r�	  j�  jg  �r�	  j  j�  �r�	  h�X   my_liner�	  �r�	  j�  j  �r�	  j�  j�  �r�	  j  j�  �r�	  hX   endr�	  �r�	  j  j�  �r�	  h�X   printr�	  �r�	  j�  j�  �r�	  j  j�  �r�	  j  j�  �r�	  j  j�  �r�	  hX   entityr�	  �r�	  j  j�  �r�	  h�X   add32csar�	  �r�	  j  j�  �r�	  hX   isr�	  �r�	  j  X
             r�	  �r�	  ji  X/   -- one stage of carry save adder for multiplierr�	  �r�	  j  j�  �r�	  j  X     r�	  �r�	  hX   portr�	  �r�	  j�  j�  �r�	  j  j�  �r�	  j  X       r�	  �r�	  h�X   br�	  �r�	  j  X          r�	  �r�	  hkj�  �r�	  j  j�  �r�	  hX   inr�	  �r�	  j  X     r�	  �r�	  hX	   std_logicr�	  �r�	  j�  j�  �r�	  j  X                         r�	  �r�	  ji  X   -- a multiplier bitr�	  �r�	  j  j�  �r�	  j  X       r�	  �r�	  h�X   ar�	  �r�	  j  X          r�	  �r�	  hkj�  �r�	  j  j�  �r�	  hX   inr�	  �r�	  j  X     r�	  �r�	  hX   std_logic_vectorr�	  �r�	  j�  j�  �r�	  j�  X   31r�	  �r�	  j  j�  �r�	  hX   downtor�	  �r�	  j  j�  �r�	  j�  j�  �r�	  j�  j  �r�	  j�  j�  �r�	  j  X     r�	  �r�	  ji  X   -- multiplicandr�	  �r�	  j  j�  �r�	  j  X       r�	  �r�	  h�X   sum_inr�	  �r 
  j  X     r
  �r
  hkj�  �r
  j  j�  �r
  hX   inr
  �r
  j  X     r
  �r
  hX   std_logic_vectorr	
  �r

  j�  j�  �r
  j�  X   31r
  �r
  j  j�  �r
  hX   downtor
  �r
  j  j�  �r
  j�  j�  �r
  j�  j  �r
  j�  j�  �r
  j  X     r
  �r
  ji  X   -- sums from previous stager
  �r
  j  j�  �r
  j  X       r
  �r
  h�X   cinr
  �r
  j  X        r
  �r
  hkj�  �r 
  j  j�  �r!
  hX   inr"
  �r#
  j  X     r$
  �r%
  hX   std_logic_vectorr&
  �r'
  j�  j�  �r(
  j�  X   31r)
  �r*
  j  j�  �r+
  hX   downtor,
  �r-
  j  j�  �r.
  j�  j�  �r/
  j�  j  �r0
  j�  j�  �r1
  j  X     r2
  �r3
  ji  X   -- carrys from previous stager4
  �r5
  j  j�  �r6
  j  X       r7
  �r8
  h�X   sum_outr9
  �r:
  j  j�  �r;
  hkj�  �r<
  j  j�  �r=
  hX   outr>
  �r?
  j  j�  �r@
  hX   std_logic_vectorrA
  �rB
  j�  j�  �rC
  j�  X   31rD
  �rE
  j  j�  �rF
  hX   downtorG
  �rH
  j  j�  �rI
  j�  j�  �rJ
  j�  j  �rK
  j�  j�  �rL
  j  X     rM
  �rN
  ji  X   -- sums to next stagerO
  �rP
  j  j�  �rQ
  j  X       rR
  �rS
  h�X   coutrT
  �rU
  j  X       rV
  �rW
  hkj�  �rX
  j  j�  �rY
  hX   outrZ
  �r[
  j  j�  �r\
  hX   std_logic_vectorr]
  �r^
  j�  j�  �r_
  j�  X   31r`
  �ra
  j  j�  �rb
  hX   downtorc
  �rd
  j  j�  �re
  j�  j�  �rf
  j�  j  �rg
  j�  j  �rh
  j�  j�  �ri
  j  j�  �rj
  ji  X   -- carrys to next stagerk
  �rl
  j  j�  �rm
  hX   endrn
  �ro
  j  j�  �rp
  h�X   add32csarq
  �rr
  j�  j�  �rs
  j  j�  �rt
  j  j�  �ru
  j  j�  �rv
  hX   ARCHITECTURErw
  �rx
  j  j�  �ry
  h�X   circuitsrz
  �r{
  j  j�  �r|
  hX   ofr}
  �r~
  j  j�  �r
  h�X   add32csar�
  �r�
  j  j�  �r�
  hX   ISr�
  �r�
  j  j�  �r�
  j  X     r�
  �r�
  hX   SIGNALr�
  �r�
  j  j�  �r�
  h�X   zeror�
  �r�
  j  j�  �r�
  hkj�  �r�
  j  j�  �r�
  hX   STD_LOGIC_VECTORr�
  �r�
  j�  j�  �r�
  j�  X   31r�
  �r�
  j  j�  �r�
  hX   downtor�
  �r�
  j  j�  �r�
  j�  j�  �r�
  j�  j  �r�
  j  j�  �r�
  hkj�  �r�
  hkj  �r�
  j  j�  �r�
  j�  X   X"00000000"r�
  �r�
  j�  j�  �r�
  j  j�  �r�
  j  X     r�
  �r�
  hX   SIGNALr�
  �r�
  j  j�  �r�
  h�X   aar�
  �r�
  j  j�  �r�
  hkj�  �r�
  j  j�  �r�
  hX   std_logic_vectorr�
  �r�
  j�  j�  �r�
  j�  X   31r�
  �r�
  j  j�  �r�
  hX   downtor�
  �r�
  j  j�  �r�
  j�  j�  �r�
  j�  j  �r�
  j  j�  �r�
  hkj�  �r�
  hkj  �r�
  j  j�  �r�
  j�  X   X"00000000"r�
  �r�
  j�  j�  �r�
  j  j�  �r�
  j  X     
  r�
  �r�
  hX	   COMPONENTr�
  �r�
  j  j�  �r�
  h�X   faddr�
  �r�
  j  X       r�
  �r�
  ji  X   -- duplicates entity portr�
  �r�
  j  j�  �r�
  j  X       r�
  �r�
  hX   PoRTr�
  �r�
  j�  j�  �r�
  h�j�	  �r�
  j  X       r�
  �r�
  hkj�  �r�
  j  j�  �r�
  hX   inr�
  �r�
  j  X     r�
  �r�
  hX	   std_logicr�
  �r�
  j�  j�  �r�
  j  j�  �r�
  j  X	            r�
  �r�
  h�j�	  �r�
  j  X       r�
  �r�
  hkj�  �r�
  j  j�  �r�
  hX   inr�
  �r�
  j  X     r�
  �r�
  hX	   std_logicr�
  �r�
  j�  j�  �r�
  j  j�  �r�
  j  X	            r�
  �r�
  h�X   cinr�
  �r�
  j  X     r�
  �r�
  hkj�  �r�
  j  j�  �r�
  hX   inr�
  �r�
  j  X     r�
  �r�
  hX	   std_logicr�
  �r�
  j�  j�  �r�
  j  j�  �r�
  j  X	            r�
  �r�
  h�X   sr�
  �r   j  X       r  �r  hkj�  �r  j  j�  �r  hX   outr  �r  j  j�  �r  hX	   std_logicr  �r	  j�  j�  �r
  j  j�  �r  j  X	            r  �r  h�X   coutr  �r  j  j�  �r  hkj�  �r  j  j�  �r  hX   outr  �r  j  j�  �r  hX	   std_logicr  �r  j�  j  �r  j�  j�  �r  j  j�  �r  j  X     r  �r  hX   endr  �r  j  j�  �r  hX	   comPonentr   �r!  j  j�  �r"  h�X   faddr#  �r$  j�  j�  �r%  j  j�  �r&  j  X     
r'  �r(  hX   beginr)  �r*  j  X     r+  �r,  ji  X   -- circuits of add32csar-  �r.  j  j�  �r/  j  X     r0  �r1  h�X   aar2  �r3  j  j�  �r4  hkj.  �r5  hkj  �r6  j  j�  �r7  h�j�	  �r8  j  j�  �r9  hX   whenr:  �r;  j  j�  �r<  h�j�	  �r=  hkj  �r>  j�  X   '1'r?  �r@  j  j�  �rA  hX   elserB  �rC  j  j�  �rD  h�X   zerorE  �rF  j  j�  �rG  hX   afterrH  �rI  j  j�  �rJ  j�  j�  �rK  j  j�  �rL  h�X   nsrM  �rN  j�  j�  �rO  j  j�  �rP  j  X     rQ  �rR  h�X   stagerS  �rT  hkj�  �rU  j  j�  �rV  hX   forrW  �rX  j  j�  �rY  h�X   IrZ  �r[  j  j�  �r\  hX   inr]  �r^  j  j�  �r_  j�  j�  �r`  j  j�  �ra  hX   torb  �rc  j  j�  �rd  j�  X   31re  �rf  j  j�  �rg  hX   generaterh  �ri  j  j�  �rj  j  X       rk  �rl  h�X   starm  �rn  hkj�  �ro  j  j�  �rp  h�X   faddrq  �rr  j  j�  �rs  hX   portrt  �ru  j  j�  �rv  hX   maprw  �rx  j�  j�  �ry  h�X   aarz  �r{  j�  j�  �r|  h�jZ  �r}  j�  j  �r~  j�  jg  �r  j  j�  �r�  h�X   sum_inr�  �r�  j�  j�  �r�  h�jZ  �r�  j�  j  �r�  j�  jg  �r�  j  j�  �r�  h�X   cinr�  �r�  j�  j�  �r�  h�jZ  �r�  j�  j  �r�  j  j�  �r�  j�  jg  �r�  j  j�  �r�  h�X   sum_outr�  �r�  j�  j�  �r�  h�jZ  �r�  j�  j  �r�  j�  jg  �r�  j  j�  �r�  h�X   coutr�  �r�  j�  j�  �r�  h�jZ  �r�  j�  j  �r�  j�  j  �r�  j�  j�  �r�  j  j�  �r�  j  X     r�  �r�  hX   endr�  �r�  j  j�  �r�  hX   generater�  �r�  j  j�  �r�  h�X   stager�  �r�  j�  j�  �r�  j  X     
r�  �r�  hX   endr�  �r�  j  j�  �r�  hX   architecturer�  �r�  j  j�  �r�  h�X   circuitsr�  �r�  j�  j�  �r�  j  j�  �r�  ji  X   -- of add32csar�  �r�  j  j�  �r�  e.