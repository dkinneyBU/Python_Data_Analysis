�]q (cpygments.token
_TokenType
qX   CommentqX   Preprocq�q�q�q}q(X   subtypesqcbuiltins
set
q	]q
�qRqX   parentqhh�q�q�q}q(hh	]q(hhhX   Multiq�q�q�q}q(hh	]q�qRqhhubhhX   Hashbangq�q�q�q}q(hh	]q �q!Rq"hhubhhX   Singleq#�q$�q%�q&}q'(hh	]q(�q)Rq*hhubhhX
   SingleLineq+�q,�q-�q.}q/(hh	]q0�q1Rq2hhubhhX   Docq3�q4�q5�q6}q7(hh	]q8�q9Rq:hhubhhX	   Directiveq;�q<�q=�q>}q?(hh	]q@�qARqBhhubhhX	   MultilineqC�qD�qE�qF}qG(hh	]qH�qIRqJhhubhhX
   SinglelineqK�qL�qM�qN}qO(hh	]qP�qQRqRhhubhhX   PreprocFileqS�qT�qU�qV}qW(hh	]qX�qYRqZhhubhhX   Specialq[�q\�q]�q^}q_(hh	]q`�qaRqbhhube�qcRqdhh)�qe�qf}qg(hh	]qh(hX   Escapeqi�qj�qk�ql}qm(hh	]qn�qoRqphhfubhX   Operatorqq�qr�qs�qt}qu(hh	]qv(hhqX   DBSqw�qx�qy�qz}q{(hh	]q|�q}Rq~hhtubhhqX   Wordq�q��q��q�}q�(hh	]q��q�Rq�hhtube�q�Rq�hhfhh�hwhzubhX   Nameq��q��q��q�}q�(hh	]q�(hh�X   Tagq��q��q��q�}q�(hh	]q��q�Rq�hh�ubhh�X   Entityq��q��q��q�}q�(hh	]q�hh�h�hw�q��q��q�}q�(hh	]q��q�Rq�hh�uba�q�Rq�hh�hwh�ubhh�X	   Exceptionq��q��q��q�}q�(hh	]q��q�Rq�hh�ubhh�X	   Decoratorq��q��q��q�}q�(hh	]q��q�Rq�hh�ubhh�X   Classq��q��q��q�}q�(hh	]q�(hh�h�hw�q��q��q�}q�(hh	]q��q�Rq�hh�ubhh�h�X   StartqÇqąqŁq�}q�(hh	]qȅq�Rq�hh�ube�q�Rq�hh�h�h�hwh�ubhh�X   Variableq͆q΅qρq�}q�(hh	]q�(hh�h�X	   AnonymousqӇqԅqՁq�}q�(hh	]q؅q�Rq�hh�ubhh�h�h��qۅq܁q�}q�(hh	]q߅q�Rq�hh�ubhh�h�X   Magicq�q�q�q�}q�(hh	]q�q�Rq�hh�ubhh�h�X   Globalq�q�q�q�}q�(hh	]q�q�Rq�hh�ubhh�h�X   Instanceq�q�q�q�}q�(hh	]q��q�Rq�hh�ube�q�Rq�hh�h�h�h�h�h�h�h�h�h�h�ubhh�X	   Attributeq��q��q��q�}r   (hh	]r  hh�h�h͇r  �r  �r  }r  (hh	]r  �r  Rr  hh�uba�r	  Rr
  hh�h�j  ubhh�X	   Namespacer  �r  �r  �r  }r  (hh	]r  �r  Rr  hh�ubhh�X   Propertyr  �r  �r  �r  }r  (hh	]r  �r  Rr  hh�ubhh�X   Symbolr  �r  �r  �r  }r  (hh	]r   �r!  Rr"  hh�ubhh�X   Classesr#  �r$  �r%  �r&  }r'  (hh	]r(  �r)  Rr*  hh�ubhh�X   Pseudor+  �r,  �r-  �r.  }r/  (hh	]r0  �r1  Rr2  hh�ubhh�X   Labelr3  �r4  �r5  �r6  }r7  (hh	]r8  �r9  Rr:  hh�ubhh�hq�r;  �r<  �r=  }r>  (hh	]r?  �r@  RrA  hh�ubhh�X   BuiltinrB  �rC  �rD  �rE  }rF  (hh	]rG  (hh�jB  j+  �rH  �rI  �rJ  }rK  (hh	]rL  �rM  RrN  hjE  ubhh�jB  X   TyperO  �rP  �rQ  �rR  }rS  (hh	]rT  �rU  RrV  hjE  ube�rW  RrX  hh�j+  jJ  jO  jR  ubhh�X   FieldrY  �rZ  �r[  �r\  }r]  (hh	]r^  �r_  Rr`  hh�ubhh�X   Otherra  �rb  �rc  �rd  }re  (hh	]rf  hh�ja  X   Memberrg  �rh  �ri  �rj  }rk  (hh	]rl  �rm  Rrn  hjd  uba�ro  Rrp  hh�jg  jj  ubhh�X   Functionrq  �rr  �rs  �rt  }ru  (hh	]rv  hh�jq  h�rw  �rx  �ry  }rz  (hh	]r{  �r|  Rr}  hjt  uba�r~  Rr  hh�h�jy  ubhh�jO  �r�  �r�  �r�  }r�  (hh	]r�  �r�  Rr�  hh�ubhh�X   Constantr�  �r�  �r�  �r�  }r�  (hh	]r�  �r�  Rr�  hh�ube�r�  Rr�  hhfh�h�jB  jE  h�h�j�  j�  h�h�h�h�h�h�jq  jt  j  j  j3  j6  j  j  ja  jd  h�h�h�h�jY  j\  j  j  j+  j.  hqj=  j#  j&  jO  j�  ubhX   Literalr�  �r�  �r�  �r�  }r�  (hh	]r�  (hj�  ja  �r�  �r�  �r�  }r�  (hh	]r�  �r�  Rr�  hj�  ubhj�  X   Charr�  �r�  �r�  �r�  }r�  (hh	]r�  �r�  Rr�  hj�  ubhj�  X   Dater�  �r�  �r�  �r�  }r�  (hh	]r�  �r�  Rr�  hj�  ubhj�  X   Scalarr�  �r�  �r�  �r�  }r�  (hh	]r�  hj�  j�  X   Plainr�  �r�  �r�  �r�  }r�  (hh	]r�  �r�  Rr�  hj�  uba�r�  Rr�  hj�  j�  j�  ubhj�  X   Stringr�  �r�  �r�  �r�  }r�  (hh	]r�  (hj�  j�  X   Interpolr�  �r�  �r�  �r�  }r�  (hh	]r�  �r�  Rr�  hj�  ubhj�  j�  X	   Delimeterr�  �r�  �r�  �r�  }r�  (hh	]r�  �r�  Rr�  hj�  ubhj�  j�  j�  �r�  �r�  �r�  }r�  (hh	]r�  �r�  Rr�  hj�  ubhj�  j�  j  �r�  �r�  �r�  }r�  (hh	]r�  �r�  Rr�  hj�  ubhj�  j�  h#�r�  �r�  �r�  }r�  (hh	]r�  �r�  Rr�  hj�  ubhj�  j�  ja  �r�  �r�  �r�  }r�  (hh	]r�  �r�  Rr�  hj�  ubhj�  j�  X   Backtickr�  �r�  �r�  �r�  }r�  (hh	]r�  �r�  Rr�  hj�  ubhj�  j�  hi�r�  �r�  �r�  }r�  (hh	]r�  �r�  Rr�  hj�  ubhj�  j�  X   Regexr�  �r   �r  �r  }r  (hh	]r  �r  Rr  hj�  ubhj�  j�  X   Momentr  �r  �r	  �r
  }r  (hh	]r  �r  Rr  hj�  ubhj�  j�  X   Booleanr  �r  �r  �r  }r  (hh	]r  �r  Rr  hj�  ubhj�  j�  X	   Characterr  �r  �r  �r  }r  (hh	]r  �r  Rr  hj�  ubhj�  j�  X	   Delimiterr  �r   �r!  �r"  }r#  (hh	]r$  �r%  Rr&  hj�  ubhj�  j�  h3�r'  �r(  �r)  }r*  (hh	]r+  �r,  Rr-  hj�  ubhj�  j�  h��r.  �r/  �r0  }r1  (hh	]r2  �r3  Rr4  hj�  ubhj�  j�  X   Affixr5  �r6  �r7  �r8  }r9  (hh	]r:  �r;  Rr<  hj�  ubhj�  j�  X   Heredocr=  �r>  �r?  �r@  }rA  (hh	]rB  �rC  RrD  hj�  ubhj�  j�  X   DoublerE  �rF  �rG  �rH  }rI  (hh	]rJ  �rK  RrL  hj�  ubhj�  j�  X   InterprM  �rN  �rO  �rP  }rQ  (hh	]rR  �rS  RrT  hj�  ubhj�  j�  X   AtomrU  �rV  �rW  �rX  }rY  (hh	]rZ  �r[  Rr\  hj�  ube�r]  Rr^  hj�  j5  j8  j�  j�  j�  j�  j  j"  h3j)  jE  jH  hij�  j=  j@  j�  j�  ja  j�  j�  j  h#j�  j  j�  j  j  j  j
  jM  jP  j  j  j�  j�  jU  jX  h�j0  ubhj�  X   Numberr_  �r`  �ra  �rb  }rc  (hh	]rd  (hj�  j_  X   Floatre  �rf  �rg  �rh  }ri  (hh	]rj  �rk  Rrl  hjb  ubhj�  j_  X   Decrm  �rn  �ro  �rp  }rq  (hh	]rr  �rs  Rrt  hjb  ubhj�  j_  X   Radixru  �rv  �rw  �rx  }ry  (hh	]rz  �r{  Rr|  hjb  ubhj�  j_  X   Octr}  �r~  �r  �r�  }r�  (hh	]r�  �r�  Rr�  hjb  ubhj�  j_  X   Binr�  �r�  �r�  �r�  }r�  (hh	]r�  �r�  Rr�  hjb  ubhj�  j_  h��r�  �r�  �r�  }r�  (hh	]r�  �r�  Rr�  hjb  ubhj�  j_  X   Hexr�  �r�  �r�  �r�  }r�  (hh	]r�  �r�  Rr�  hjb  ubhj�  j_  X   Integerr�  �r�  �r�  �r�  }r�  (hh	]r�  h(j�  j_  j�  X   Longr�  tr�  �r�  �r�  }r�  (hh	]r�  �r�  Rr�  hj�  uba�r�  Rr�  hjb  j�  j�  ubhj�  j_  X   Decimalr�  �r�  �r�  �r�  }r�  (hh	]r�  �r�  Rr�  hjb  ube�r�  Rr�  hj�  j�  j�  je  jh  j�  j�  j�  j�  j}  j�  ju  jx  h�j�  j�  j�  jm  jp  ube�r�  Rr�  hhfj�  j�  j_  jb  j�  j�  j�  j�  ja  j�  j�  j�  ubhX   Genericr�  �r�  �r�  �r�  }r�  (hh	]r�  (hj�  X   Errorr�  �r�  �r�  �r�  }r�  (hh	]r�  �r�  Rr�  hj�  ubhj�  X
   Subheadingr�  �r�  �r�  �r�  }r�  (hh	]r�  �r�  Rr�  hj�  ubhj�  X	   Tracebackr�  �r�  �r�  �r�  }r�  (hh	]r�  �r�  Rr�  hj�  ubhj�  X   Outputr�  �r�  �r�  �r�  }r�  (hh	]r�  �r�  Rr�  hj�  ubhj�  X   Promptr�  �r�  �r�  �r�  }r�  (hh	]r�  �r�  Rr�  hj�  ubhj�  X   Deletedr�  �r�  �r�  �r�  }r�  (hh	]r�  �r�  Rr�  hj�  ubhj�  X   Insertedr�  �r�  �r�  �r�  }r�  (hh	]r�  �r�  Rr�  hj�  ubhj�  X   Headingr�  �r�  �r�  �r�  }r�  (hh	]r�  �r�  Rr�  hj�  ubhj�  X   Strongr�  �r�  �r   �r  }r  (hh	]r  �r  Rr  hj�  ubhj�  X   Emphr  �r  �r  �r	  }r
  (hh	]r  �r  Rr  hj�  ube�r  Rr  hhfj�  j�  j  j	  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j�  j  j�  j�  j�  j�  ubhj�  �r  �r  �r  }r  (hh	]r  �r  Rr  hhfubhX   Keywordr  �r  �r  �r  }r  (hh	]r  (hj  h�r  �r  �r  }r   (hh	]r!  �r"  Rr#  hj  ubhj  j  �r$  �r%  �r&  }r'  (hh	]r(  �r)  Rr*  hj  ubhj  jO  �r+  �r,  �r-  }r.  (hh	]r/  �r0  Rr1  hj  ubhj  X   PreProcr2  �r3  �r4  �r5  }r6  (hh	]r7  �r8  Rr9  hj  ubhj  X   Controlr:  �r;  �r<  �r=  }r>  (hh	]r?  �r@  RrA  hj  ubhj  j�  �rB  �rC  �rD  }rE  (hh	]rF  �rG  RrH  hj  ubhj  j  �rI  �rJ  �rK  }rL  (hh	]rM  �rN  RrO  hj  ubhj  j+  �rP  �rQ  �rR  }rS  (hh	]rT  �rU  RrV  hj  ubhj  X   DeclarationrW  �rX  �rY  �rZ  }r[  (hh	]r\  �r]  Rr^  hj  ubhj  X   Reservedr_  �r`  �ra  �rb  }rc  (hh	]rd  �re  Rrf  hj  ube�rg  Rrh  hhfj�  jD  jW  jZ  j  jK  j+  jR  j_  jb  jO  j-  j:  j=  j  j&  j2  j5  hj  ubhja  �ri  �rj  �rk  }rl  (hh	]rm  �rn  Rro  hhfubhX   Textrp  �rq  �rr  �rs  }rt  (hh	]ru  (hjp  X   Rootrv  �rw  �rx  �ry  }rz  (hh	]r{  �r|  Rr}  hjs  ubhjp  j  �r~  �r  �r�  }r�  (hh	]r�  �r�  Rr�  hjs  ubhjp  X   Ragr�  �r�  �r�  �r�  }r�  (hh	]r�  �r�  Rr�  hjs  ubhjp  X
   Whitespacer�  �r�  �r�  �r�  }r�  (hh	]r�  �r�  Rr�  hjs  ubhjp  X   Beerr�  �r�  �r�  �r�  }r�  (hh	]r�  �r�  Rr�  hjs  ubhjp  X   Punctuationr�  �r�  �r�  �r�  }r�  (hh	]r�  �r�  Rr�  hjs  ube�r�  Rr�  hhfj�  j�  j  j�  j�  j�  jv  jy  j�  j�  j�  j�  ubhhj�  �r�  �r�  �r�  }r�  (hh	]r�  hj�  X	   Indicatorr�  �r�  �r�  �r�  }r�  (hh	]r�  �r�  Rr�  hj�  uba�r�  Rr�  hhfj�  j�  ube�r�  Rr�  jp  js  hihlj�  j  ja  jk  j  j  h�h�j�  j�  j�  j�  hqhthhj�  j�  X   Tokenr�  hfj�  j�  j_  jb  ubhhhChFhhhShVh#h&h[h^h;h>h+h.h3h6hhhKhNububX   #ifdef ARCH_ARM
r�  �r�  j  X   archr�  �r�  js  X    r�  �r�  j  X   arm11r�  �r�  js  X   
r�  �r�  hX   #else
r�  �r�  j  X   archr�  �r�  js  j�  �r�  j  X   ia32r�  �r�  js  j�  �r�  hX   #endif
r�  �r�  js  j�  �r�  j  X   objectsr�  �r�  js  j�  �r�  j�  X   {r�  �r�  js  X   
  r�  �r�  h�X   my_epr�  �r�  js  j�  �r�  j�  X   =r�  �r�  js  j�  �r�  j-  X   epr�  �r�  js  j�  �r�  hX   /* A synchronous endpoint */r�  �r�  js  X   

  r�  �r�  hX   /* Two thread control blocks */r�  �r�  js  X   
  r�  �r�  h�X   tcb1r�  �r�  js  j�  �r�  j�  j�  �r�  js  j�  �r�  j-  X   tcbr�  �r�  js  X   
  r�  �r�  h�X   tcb2r�  �r�  js  j�  �r�  j�  j�  �r�  js  j�  �r�  j-  X   tcbr�  �r�  js  X   

  r�  �r�  hX$   /* Four frames of physical memory */r�  �r�  js  X   
  r�  �r�  h�X   frame1r�  �r�  js  j�  �r�  j�  j�  �r�  js  j�  �r   j-  X   framer  �r  js  j�  �r  j�  X   (r  �r  jb  X   4kr  �r  j�  X   )r  �r	  js  X   
  r
  �r  h�X   frame2r  �r  js  j�  �r  j�  j�  �r  js  j�  �r  j-  X   framer  �r  js  j�  �r  j�  j  �r  jb  X   4kr  �r  j�  j  �r  js  X   
  r  �r  h�X   frame3r  �r  js  j�  �r  j�  j�  �r  js  j�  �r  j-  X   framer  �r   js  j�  �r!  j�  j  �r"  jb  X   4kr#  �r$  j�  j  �r%  js  X   
  r&  �r'  h�X   frame4r(  �r)  js  j�  �r*  j�  j�  �r+  js  j�  �r,  j-  X   framer-  �r.  js  j�  �r/  j�  j  �r0  jb  X   4kr1  �r2  j�  j  �r3  js  X   

  r4  �r5  hX   /* Two page tables */r6  �r7  js  X   
  r8  �r9  h�X   pt1r:  �r;  js  j�  �r<  j�  j�  �r=  js  j�  �r>  j-  X   ptr?  �r@  js  X   
  rA  �rB  h�X   pt2rC  �rD  js  j�  �rE  j�  j�  �rF  js  j�  �rG  j-  X   ptrH  �rI  js  X   

  rJ  �rK  hX   /* Two page directories */rL  �rM  js  X   
  rN  �rO  h�X   pd1rP  �rQ  js  j�  �rR  j�  j�  �rS  js  j�  �rT  j-  X   pdrU  �rV  js  X   
  rW  �rX  h�X   pd2rY  �rZ  js  j�  �r[  j�  j�  �r\  js  j�  �r]  j-  X   pdr^  �r_  js  X   

  r`  �ra  hX   /* Two capability nodes */rb  �rc  js  X   
  rd  �re  h�X   cnode1rf  �rg  js  j�  �rh  j�  j�  �ri  js  j�  �rj  j-  X   cnoderk  �rl  js  j�  �rm  j�  j  �rn  jb  X   2ro  �rp  js  j�  �rq  jb  X   bitsrr  �rs  j�  j  �rt  js  X   
  ru  �rv  h�X   cnode2rw  �rx  js  j�  �ry  j�  j�  �rz  js  j�  �r{  j-  X   cnoder|  �r}  js  j�  �r~  j�  j  �r  jb  X   3r�  �r�  js  j�  �r�  jb  X   bitsr�  �r�  j�  j  �r�  js  j�  �r�  j�  X   }r�  �r�  js  j�  �r�  j  X   capsr�  �r�  js  j�  �r�  j�  j�  �r�  js  X   
  r�  �r�  h�X   cnode1r�  �r�  js  j�  �r�  j�  j�  �r�  js  X   
    r�  �r�  j�  X   0x1r�  �r�  j�  X   :r�  �r�  js  j�  �r�  h�X   frame1r�  �r�  js  j�  �r�  j�  j  �r�  jb  X   RWr�  �r�  j�  j  �r�  js  j�  �r�  hX   /* read/write */r�  �r�  js  X   
    r�  �r�  j�  X   0x2r�  �r�  j�  j�  �r�  js  j�  �r�  h�X   my_epr�  �r�  js  j�  �r�  j�  j  �r�  jb  X   Rr�  �r�  j�  j  �r�  js  X      r�  �r�  hX   /* read-only */r�  �r�  js  X   
  r�  �r�  j�  j�  �r�  js  X   
  r�  �r�  h�X   cnode2r�  �r�  js  j�  �r�  j�  j�  �r�  js  X   
    r�  �r�  j�  X   0x1r�  �r�  j�  j�  �r�  js  j�  �r�  h�X   my_epr�  �r�  js  j�  �r�  j�  j  �r�  jb  X   Wr�  �r�  j�  j  �r�  js  X      r�  �r�  hX   /* write-only */r�  �r�  js  X   
  r�  �r�  j�  j�  �r�  js  X   
  r�  �r�  h�X   tcb1r�  �r�  js  j�  �r�  j�  j�  �r�  js  X   
    r�  �r�  jb  X   vspacer�  �r�  j�  j�  �r�  js  j�  �r�  h�X   pd1r�  �r�  js  X   
    r�  �r�  jb  X   ipc_buffer_slotr�  �r�  j�  j�  �r�  js  j�  �r�  h�X   frame1r�  �r�  js  X   
    r�  �r�  jb  X   cspacer�  �r�  j�  j�  �r�  js  j�  �r�  h�X   cnode1r�  �r�  js  X   
  r�  �r�  j�  j�  �r�  js  X   
  r�  �r�  h�X   pd1r�  �r�  js  j�  �r�  j�  j�  �r�  js  X   
    r�  �r�  j�  X   0x10r�  �r�  j�  j�  �r�  js  j�  �r�  h�X   pt1r   �r  js  X   
  r  �r  j�  j�  �r  js  X   
  r  �r  h�X   pt1r  �r  js  j�  �r	  j�  j�  �r
  js  X   
    r  �r  j�  X   0x8r  �r  j�  j�  �r  js  j�  �r  h�X   frame1r  �r  js  j�  �r  j�  j  �r  jb  X   RWr  �r  j�  j  �r  js  X   
    r  �r  j�  X   0x9r  �r  j�  j�  �r  js  j�  �r  h�X   frame2r  �r  js  j�  �r   j�  j  �r!  jb  j�  �r"  j�  j  �r#  js  X   
  r$  �r%  j�  j�  �r&  js  X   
  r'  �r(  h�X   tcb2r)  �r*  js  j�  �r+  j�  j�  �r,  js  X   
    r-  �r.  jb  X   vspacer/  �r0  j�  j�  �r1  js  j�  �r2  h�X   pd2r3  �r4  js  X   
    r5  �r6  jb  X   ipc_buffer_slotr7  �r8  j�  j�  �r9  js  j�  �r:  h�X   frame3r;  �r<  js  X   
    r=  �r>  jb  X   cspacer?  �r@  j�  j�  �rA  js  j�  �rB  h�X   cnode2rC  �rD  js  X   
  rE  �rF  j�  j�  �rG  js  X   
  rH  �rI  h�X   pd2rJ  �rK  js  j�  �rL  j�  j�  �rM  js  X   
    rN  �rO  j�  X   0x10rP  �rQ  j�  j�  �rR  js  j�  �rS  h�X   pt2rT  �rU  js  X   
  rV  �rW  j�  j�  �rX  js  X   
  rY  �rZ  h�X   pt2r[  �r\  js  j�  �r]  j�  j�  �r^  js  X   
    r_  �r`  j�  X   0x10ra  �rb  j�  j�  �rc  js  j�  �rd  h�X   frame3re  �rf  js  j�  �rg  j�  j  �rh  jb  X   RWri  �rj  j�  j  �rk  js  X   
    rl  �rm  j�  X   0x12rn  �ro  j�  j�  �rp  js  j�  �rq  h�X   frame4rr  �rs  js  j�  �rt  j�  j  �ru  jb  j�  �rv  j�  j  �rw  js  X   
  rx  �ry  j�  j�  �rz  js  j�  �r{  j�  j�  �r|  js  j�  �r}  e.